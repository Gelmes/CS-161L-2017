`timescale 1ns / 1ps

module CAMArray(
    );


endmodule
